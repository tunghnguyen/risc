module inst_mem (
    input wire [31:0] addr,
    input wire clk,
    output reg [31:0] inst
);



endmodule
