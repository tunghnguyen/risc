module dat_mem (
    input wire [31:0] addr,
    input wire [31:0] w_dat,
    input wire mem_read,
    input wire mem_write,
    input wire clk,
    output reg [31:0] r_dat
);



endmodule
