module risc ();

endmodule
