module risc;

endmodule
